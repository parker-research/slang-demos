module m;
struct {
    int i;
    logic l;
} s;
endmodule
